// ��Ʈ ������
// ���� ���� �ð��� ���� �Ǻ� ������ ���� ��ȣ ����

module note_gen (
    input clk,
    input rst,
    input [31:0] i_cur_time, // game_timer���� ���� ���� �ð� (ms)
    
    output reg o_note_t1,    // Track 1 (����) ��Ʈ ���� ��ȣ (1ƽ ���� 1)
    output reg o_note_t2,    // Track 2 (�Ʒ���) ��Ʈ ���� ��ȣ
    output reg o_game_end    // �뷡�� �������� �˸��� ��ȣ
);

    // ==========================================
    // �Ǻ� ������ �ϵ��ڵ�
    // ==========================================
    // ��Ʈ ����
    parameter NOTE_COUNT = 10;
    
    reg [31:0] note_time [0:NOTE_COUNT-1]; // �ð� ����
    reg [1:0]  note_track [0:NOTE_COUNT-1]; // Ʈ�� ���� (1:����, 2:�Ʒ���, 3:����)

    initial begin
        // {�ð�(ms), Ʈ��}
        // LCD ������ ������ ���� ���������� ���µ� �ɸ��� �ð��� ����ؼ� ��ġ
        // ��: ��ũ�� �ӵ��� �����ٸ�, �����ϰ� ���� �ð����� ���� ���� �����ؾ� ��
        
        // �ϴ��� '���� �ð�' �������� �ۼ��� ���ô�.
        note_time[0] = 1000; note_track[0] = 1; // 1��: ����
        note_time[1] = 2000; note_track[1] = 2; // 2��: �Ʒ���
        note_time[2] = 2500; note_track[2] = 1; 
        note_time[3] = 3000; note_track[3] = 2;
        note_time[4] = 3500; note_track[4] = 1;
        note_time[5] = 4000; note_track[5] = 3; // 4��: ���� ġ��!
        note_time[6] = 5000; note_track[6] = 1;
        note_time[7] = 5500; note_track[7] = 2;
        note_time[8] = 6000; note_track[8] = 1;
        note_time[9] = 7000; note_track[9] = 3; // ������ ���� ġ��
    end

    // ==========================================
    // ������ ���� (FSM)
    // ==========================================
    reg [31:0] note_idx; // ���� �� ��° ��Ʈ�� ��ٸ��� ������ (������)

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            note_idx <= 0;
            o_note_t1 <= 0;
            o_note_t2 <= 0;
            o_game_end <= 0;
        end else begin
            o_note_t1 <= 0;
            o_note_t2 <= 0;

            // �뷡�� ���� �� �����ٸ�
            if (note_idx < NOTE_COUNT) begin
                // ���� �ð��� ��Ʈ�� �ð��� ���ų� ��������? (������ ��� ��� >= ���)
                if (i_cur_time >= note_time[note_idx]) begin
                    
                    // �ش� Ʈ���� ��ȣ �߻�
                    if (note_track[note_idx] == 1 || note_track[note_idx] == 3) 
                        o_note_t1 <= 1;
                    
                    if (note_track[note_idx] == 2 || note_track[note_idx] == 3) 
                        o_note_t2 <= 1;

                    // ���� ��Ʈ�� ������ �̵�
                    note_idx <= note_idx + 1;
                end
            end else begin
                // ��� ��Ʈ�� �� �������� ���� ���� ��ȣ
                // (������ ��Ʈ ������ ���� �ڿ� ������ ������ ���⼭ �ð� üũ�� �� �ص� ��)
                o_game_end <= 1;
            end
        end
    end

endmodule