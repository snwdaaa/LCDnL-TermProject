module u_game_7_segment (
    input clk,              // �ý��� Ŭ��
    input rst,              // ����
    input [1:0] i_judge,    // ���� �Է� (00:None, 01:Miss, 10:Normal, 11:Perfect)
    
    output reg [7:0] o_seg, // 7-Segment ������ �� (a,b,c,d,e,f,g,dp)
    output reg [7:0] o_com  // 7-Segment �ڸ��� ���� �� (Common)
);

    // ====================================================
    // Part 1: ���� ��� ���� (Score Logic)
    // ====================================================
    reg [13:0] score;       // ���� ���� ���� �������� (0 ~ 9999)
    reg [1:0] prev_judge;   // Edge Detection�� ���� ���� ����

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            score <= 0;
            prev_judge <= 0;
        end else begin
            // [Edge Detection] ���� ��ȣ�� ���ϴ� ����(Rising Edge)�� ����
            if (i_judge != 0 && i_judge != prev_judge) begin
                case (i_judge)
                    2'b11: score <= score + 2; // Perfect: +2��
                    2'b10: score <= score + 1; // Normal: +1��
                    2'b01: score <= score;     // Miss: 0�� (�״��)
                    default: score <= score;
                endcase
            end
            prev_judge <= i_judge; // ���� ���¸� ���ŷ� ����
        end
    end

    // ====================================================
    // Part 2: 10���� �и� (Binary to BCD)
    // ====================================================
    // 4�ڸ� ���� �и� (��: 1234 -> 1, 2, 3, 4)
    wire [3:0] digit_1 = score % 10;
    wire [3:0] digit_10 = (score / 10) % 10;
    wire [3:0] digit_100 = (score / 100) % 10;
    wire [3:0] digit_1000 = (score / 1000) % 10;

    // ====================================================
    // Part 3: ��ĳ�� �� ���÷��� ���� (Display Driver)
    // ====================================================
    reg [16:0] scan_cnt; // ��ĵ �ӵ� ������ Ÿ�̸�
    
    always @(posedge clk or posedge rst) begin
        if (rst) scan_cnt <= 0;
        else scan_cnt <= scan_cnt + 1;
    end

    // Ÿ�̸��� ���� 2��Ʈ�� ����Ͽ� 00->01->10->11 ������ �ڸ��� ��ȸ
    wire [1:0] scan_idx = scan_cnt[16:15];
    reg [3:0] current_digit_value; // ���� ���� �ڸ��� ǥ���� ����

    // 1. �ڸ��� ���� (Active Low ����: 0�� �� ����)
    always @(*) begin
        // �ϴ� �� ���� ���� (�ʱ�ȭ)
        o_com = 8'b11111111; 
        
        case (scan_idx)
            2'b00: begin
                o_com = 8'b11111110;       // ù ��° �ڸ� (���� �ڸ�, ����)
                current_digit_value = digit_1;
            end
            2'b01: begin
                o_com = 8'b11111101;       // �� ��° �ڸ� (���� �ڸ�)
                current_digit_value = digit_10;
            end
            2'b10: begin
                o_com = 8'b11111011;       // �� ��° �ڸ� (���� �ڸ�)
                current_digit_value = digit_100;
            end
            2'b11: begin
                o_com = 8'b11110111;       // �� ��° �ڸ� (õ�� �ڸ�, ����)
                current_digit_value = digit_1000;
            end
        endcase
    end

    // 2. ���� ���� ���ڵ� (Active Low ����: 0�� �� ����)
    // a~g, dp ����
    always @(*) begin
        case (current_digit_value)
            4'h0: o_seg = 8'b11000000; // 0
            4'h1: o_seg = 8'b11111001; // 1
            4'h2: o_seg = 8'b10100100; // 2
            4'h3: o_seg = 8'b10110000; // 3
            4'h4: o_seg = 8'b10011001; // 4
            4'h5: o_seg = 8'b10010010; // 5
            4'h6: o_seg = 8'b10000010; // 6
            4'h7: o_seg = 8'b11111000; // 7
            4'h8: o_seg = 8'b10000000; // 8
            4'h9: o_seg = 8'b10010000; // 9
            default: o_seg = 8'b11111111; // Off
        endcase
    end

endmodule