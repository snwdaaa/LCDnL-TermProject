module lcd_ctrl (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,              // ����
    input i_tick,           // 1ms ƽ (��ũ�� �ӵ� ������)
    
    // ��Ʈ ���� ��ȣ (from note_gen)
    input i_note_t1,        // ���� (Track 1) ��Ʈ
    input i_note_t2,        // �Ʒ��� (Track 2) ��Ʈ
    
    input [31:0] i_gen_pitch, // note_gen���� ���� ����
    
    // [NEW] ���� ���� �� ��Ʈ�� ����� ���� �Է� ��ȣ
    input i_clear_t1_perf, // Track 1 Perfect ��ġ(0��) ������
    input i_clear_t1_norm, // Track 1 Normal ��ġ(1��) ������
    input i_clear_t2_perf,
    input i_clear_t2_norm,
    
    // ���� ���� ��ȣ
    input i_game_start, // 0: ��� ȭ��, 1: ���� ����
    input i_game_over,  // 0: ���� ��, 1: ���� ����
    
    // LCD �ϵ���� �� (���� �ɿ� ����)
    output reg o_lcd_rs,    // 0:���, 1:������
    output reg o_lcd_rw,    // 0:����, 1:�б� (�׻� 0)
    output reg o_lcd_e,     // Enable �޽�
    output reg [7:0] o_lcd_data, // ������ ����
    
    // [NEW] ���� ���� ���� �˸� ��ȣ
    output o_hit_t1,      // [0�� ĭ] Perfect �� ����
    output o_pre_hit_t1,  // [1�� ĭ] Normal �� ����
    output o_hit_t2,      
    output o_pre_hit_t2,  
    
    // [NEW] ��ħ(Miss) �˸� ��ȣ
    output reg o_miss_t1, 
    output reg o_miss_t2,
    
    // ���� �������� �ִ� ��Ʈ�� ���� ��
    output reg [31:0] o_curr_pitch_t1, 
    output reg [31:0] o_curr_pitch_t2
);

    // ====================================================
    // [Part 1] ��Ʈ ��ũ�Ѹ� �� ���� ���� ����
    // ====================================================
    
    // 1. ȭ�� ���� (16ĭ x 2��)
    reg [7:0] line1 [0:15]; // ����
    reg [7:0] line2 [0:15]; // �Ʒ���
    
    // ���� ����
    reg [31:0] pitch_buf_t1 [0:15];
    reg [31:0] pitch_buf_t2 [0:15];

    // 2. ��Ʈ ĸó (Note Capture)
    reg r_catch_t1, r_catch_t2;
    reg [31:0] r_catch_pitch;

    // 3. ��ũ�� Ÿ�̸� (Scroll Timer)
    parameter SCROLL_SPEED = 300; 
    reg [31:0] scroll_cnt;
    wire scroll_en;

    always @(posedge clk or posedge rst) begin
        if (rst) scroll_cnt <= 0;
        else if (i_tick) begin
            if (scroll_cnt >= SCROLL_SPEED - 1) scroll_cnt <= 0;
            else scroll_cnt <= scroll_cnt + 1;
        end
    end
    assign scroll_en = (i_tick && (scroll_cnt == 0));

    // 4. ���� ������Ʈ (�ٽ� ����: �̵�, Miss, Clear)
    integer i;
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            // ���� �� "Press Start..." ������ �ʱ�ȭ
            // "Press Start Btn " (16����)
            line1[0]<="P"; line1[1]<="r"; line1[2]<="e"; line1[3]<="s"; 
            line1[4]<="s"; line1[5]<=" "; line1[6]<="S"; line1[7]<="t"; 
            line1[8]<="a"; line1[9]<="r"; line1[10]<="t"; line1[11]<=" "; 
            line1[12]<="B"; line1[13]<="t"; line1[14]<="n"; line1[15]<=" ";
            
            // �ʱ�ȭ
            for (i=0; i<16; i=i+1) begin
                line2[i] <= 8'h20; // �Ʒ��� ����    
                pitch_buf_t1[i] <= 0; pitch_buf_t2[i] <= 0;
            end
            r_catch_t1 <= 0; r_catch_t2 <= 0; r_catch_pitch <= 0;
            o_miss_t1 <= 0; o_miss_t2 <= 0;
        end
        else begin
            // (1) �켱���� 1: ���� ���� ȭ��
            if (i_game_over) begin
                // "   Game Over!   "
                line1[0]<=" "; line1[1]<=" "; line1[2]<=" "; line1[3]<="G"; 
                line1[4]<="a"; line1[5]<="m"; line1[6]<="e"; line1[7]<=" "; 
                line1[8]<="O"; line1[9]<="v"; line1[10]<="e"; line1[11]<="r"; 
                line1[12]<="!"; line1[13]<=" "; line1[14]<=" "; line1[15]<=" ";
                
                for (i=0; i<16; i=i+1) begin
                    line2[i] <= 8'h20; // �Ʒ��� ���� 
                end
            end
            // (2) �켱���� 2: ���� ��� ȭ�� (���� ��)
            else if (i_game_start == 0) begin
                // ���°� �����ϰ� "Press Start Btn " ����
                line1[0]<="P"; line1[1]<="r"; line1[2]<="e"; line1[3]<="s"; 
                line1[4]<="s"; line1[5]<=" "; line1[6]<="S"; line1[7]<="t"; 
                line1[8]<="a"; line1[9]<="r"; line1[10]<="t"; line1[11]<=" "; 
                line1[12]<="B"; line1[13]<="t"; line1[14]<="n"; line1[15]<=" ";
            end        
            // (3) �켱���� 3: ���� �÷��� (���� ��ũ�� ����)
            
            else begin
                // (1) Miss ���� �÷��� �ʱ�ȭ (�� Ŭ������ ����)
                o_miss_t1 <= 0; 
                o_miss_t2 <= 0;
    
                // (2) ��ũ�� ���� (Shift)
                if (scroll_en) begin
                    // �̵��ϱ� ���� �� ��(0��)�� ��Ʈ�� �־����� -> Miss �߻�!
                    if (line1[0] == 8'h4F) o_miss_t1 <= 1;
                    if (line2[0] == 8'h4F) o_miss_t2 <= 1;
    
                    // [�������� �̵�]
                    for (i=0; i<15; i=i+1) begin
                        line1[i] <= line1[i+1];
                        line2[i] <= line2[i+1];
                        pitch_buf_t1[i] <= pitch_buf_t1[i+1];
                        pitch_buf_t2[i] <= pitch_buf_t2[i+1];
                    end
                    
                    // [������ �� ä���]
                    line1[15] <= (r_catch_t1) ? 8'h4F : 8'h20;
                    line2[15] <= (r_catch_t2) ? 8'h4F : 8'h20;
                    pitch_buf_t1[15] <= (r_catch_t1) ? r_catch_pitch : 0;
                    pitch_buf_t2[15] <= (r_catch_t2) ? r_catch_pitch : 0;
                    
                    // ĸó �ʱ�ȭ
                    r_catch_t1 <= 0; r_catch_t2 <= 0;
                end 
                else begin
                    // ��ũ���� �ƴ� ��: �� ��Ʈ ĸó
                    if (i_note_t1) begin r_catch_t1 <= 1; r_catch_pitch <= i_gen_pitch; end
                    if (i_note_t2) begin r_catch_t2 <= 1; r_catch_pitch <= i_gen_pitch; end
                end
    
                // (3) [NEW] ��Ʈ ����� (Clear Note) - ���� ���� �� ����
                // Judgement ��⿡�� ��û�� ���� �ش� ĭ�� �������� ���
                
                // Track 1 Clear
                if (i_clear_t1_perf) begin line1[0] <= 8'h20; pitch_buf_t1[0] <= 0; end
                if (i_clear_t1_norm) begin line1[1] <= 8'h20; pitch_buf_t1[1] <= 0; end
                
                // Track 2 Clear
                if (i_clear_t2_perf) begin line2[0] <= 8'h20; pitch_buf_t2[0] <= 0; end
                if (i_clear_t2_norm) begin line2[1] <= 8'h20; pitch_buf_t2[1] <= 0; end
            end
        end
    end
    
    // ====================================================
    // [Part 3] ���� ���� ��ȣ ���
    // ====================================================
    // 'O' (0x4F) ���ڰ� �ִ��� Ȯ��
    assign o_hit_t1     = (line1[0] == 8'h4F); // 0�� ĭ (Perfect)
    assign o_pre_hit_t1 = (line1[1] == 8'h4F); // 1�� ĭ (Normal)
    
    assign o_hit_t2     = (line2[0] == 8'h4F);
    assign o_pre_hit_t2 = (line2[1] == 8'h4F);
    
    // ���� ��� ����: Perfect(0��) �Ǵ� Normal(1��) ��ġ�� ���� ���� ����
    always @(*) begin
        // [Track 1]
        if (pitch_buf_t1[0] > 0)       
            o_curr_pitch_t1 = pitch_buf_t1[0]; // 0���� ��Ʈ�� ������ 1���� (Perfect)
        else if (pitch_buf_t1[1] > 0)  
            o_curr_pitch_t1 = pitch_buf_t1[1]; // 1���� ��Ʈ�� ������ 2���� (Normal)
        else                           
            o_curr_pitch_t1 = 0;               // �� �� ������ 0

        // [Track 2]
        if (pitch_buf_t2[0] > 0)       
            o_curr_pitch_t2 = pitch_buf_t2[0];
        else if (pitch_buf_t2[1] > 0)  
            o_curr_pitch_t2 = pitch_buf_t2[1];
        else                           
            o_curr_pitch_t2 = 0;
    end

    // ====================================================
    // [Part 2] LCD ����̹� (Hardware Control FSM) - ���� ����
    // ====================================================
    
    // ���� ����
    localparam S_INIT       = 0;
    localparam S_CMD_PRE    = 1;
    localparam S_CMD_SEND   = 2;
    localparam S_CMD_HOLD   = 3;
    localparam S_DATA_PRE   = 4;
    localparam S_DATA_SEND  = 5;
    localparam S_DATA_HOLD  = 6;
    
    reg [3:0] state;
    reg [4:0] init_step;
    reg [4:0] char_idx;
    reg [31:0] delay_cnt;
    
    parameter DLY_2MS = 100000;
    parameter DLY_50US = 2500;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= S_INIT;
            init_step <= 0;
            char_idx <= 0;
            delay_cnt <= 0;
            o_lcd_e <= 0;
            o_lcd_rs <= 0;
            o_lcd_rw <= 0;
            o_lcd_data <= 0;
        end else begin
            case (state)
                S_INIT: begin
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > DLY_2MS * 10) begin 
                        delay_cnt <= 0;
                        state <= S_CMD_PRE;
                    end
                end

                S_CMD_PRE: begin
                    o_lcd_rs <= 0; 
                    o_lcd_rw <= 0; 
                    o_lcd_e  <= 0;
                    case (init_step)
                        0: o_lcd_data <= 8'h38;
                        1: o_lcd_data <= 8'h0C;
                        2: o_lcd_data <= 8'h06;
                        3: o_lcd_data <= 8'h01;
                        4: o_lcd_data <= 8'h80;
                        5: o_lcd_data <= 8'hC0;
                        default: o_lcd_data <= 8'h80;
                    endcase
                    state <= S_CMD_SEND;
                end

                S_CMD_SEND: begin
                    o_lcd_e <= 1;
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > 50) begin 
                        delay_cnt <= 0;
                        state <= S_CMD_HOLD;
                    end
                end
                
                S_CMD_HOLD: begin
                    o_lcd_e <= 0;
                    delay_cnt <= delay_cnt + 1;
                    if ((init_step == 3 && delay_cnt > DLY_2MS) || 
                        (init_step != 3 && delay_cnt > DLY_50US)) begin
                        delay_cnt <= 0;
                        if (init_step < 4) begin
                            init_step <= init_step + 1;
                            state <= S_CMD_PRE;
                        end else begin
                            if (init_step == 4) begin
                                char_idx <= 0;
                                state <= S_DATA_PRE; 
                            end else if (init_step == 5) begin
                                char_idx <= 16;
                                state <= S_DATA_PRE;
                            end
                        end
                    end
                end

                S_DATA_PRE: begin
                    o_lcd_rs <= 1; 
                    o_lcd_rw <= 0;
                    o_lcd_e  <= 0;
                    if (char_idx < 16) 
                        o_lcd_data <= line1[char_idx];
                    else 
                        o_lcd_data <= line2[char_idx - 16];
                    state <= S_DATA_SEND;
                end

                S_DATA_SEND: begin
                    o_lcd_e <= 1;
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > 50) begin
                        delay_cnt <= 0;
                        state <= S_DATA_HOLD;
                    end
                end

                S_DATA_HOLD: begin
                    o_lcd_e <= 0;
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > DLY_50US) begin
                        delay_cnt <= 0;
                        if (char_idx == 15) begin
                            init_step <= 5; 
                            state <= S_CMD_PRE;
                        end else if (char_idx == 31) begin
                            init_step <= 4; 
                            state <= S_CMD_PRE;
                        end else begin
                            char_idx <= char_idx + 1;
                            state <= S_DATA_PRE;
                        end
                    end
                end
            endcase
        end
    end

endmodule