module sys_base (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,              // ����
    
    // �ǿ��� ���� ��� (������ ���� �ǵ��)
    output o_piezo,
    
    // LCD ���� ��
    output o_lcd_rs,
    output o_lcd_rw,
    output o_lcd_e,
    output [7:0] o_lcd_data,
    
    // Ǯ�÷� LED ��� ��Ʈ
    output [3:0] o_fcl_r, 
    output [3:0] o_fcl_g, 
    output [3:0] o_fcl_b,
    
    // ���� 7-Segment�� ��� �� (Single)
    output [7:0] o_single_seg, 

    // 8-Array Segment�� ��� �� (Array)
    output [7:0] o_array_seg, // a~g, dp ����
    output [7:0] o_array_com, // Digit Select
    
    // ��ư �Է�
    input [3:0] i_btn       // ��ư �Է� 4��
);

    // ====================================================
    // 1. ���� ��ȣ ����
    // ====================================================
    wire w_game_tick;       // 1ms ƽ
    wire [31:0] w_cur_time; // ���� ���� �ð�
    
    // ��Ʈ ��ȣ
    wire w_note_t1;         // ���� ��Ʈ
    wire w_note_t2;         // �Ʒ��� ��Ʈ
    wire w_game_end;
    
    // ��ư ��ȣ (ä�͸� ���ŵ�)
    wire w_start_btn;
    wire w_restart_btn;
    wire [1:0] w_play_btn;  // [1]: Down(Track2), [0]: Up(Track1)
    
    // �ǿ��� ���� ��ȣ (Judgement -> Piezo)
    wire w_play_en;         // �Ҹ� ��� Enable
    wire [31:0] w_cnt_limit;// ����� ���ļ� ��
    
    // ���� ��� ��ȣ (���� ��� �� ��, ���� Ȯ���)
    wire [1:0] w_judge;     
    
    // LCD ������ ���� ��ȣ
    wire w_hit_t1, w_hit_t2;
    
    wire [31:0] w_gen_pitch;        // note_gen -> lcd_ctrl
    wire [31:0] w_curr_pitch_t1;    // lcd_ctrl -> logic
    wire [31:0] w_curr_pitch_t2;    // lcd_ctrl -> logic
    
    // ��� �� ������ ���� ��ȣ�� (Wire)
    wire [1:0] w_judge;         // ���� ��� (Judge -> Score, LED)
    wire [1:0] w_judge_hold;
    wire [15:0] w_total_score;  // ���� ���� (Score -> 7-Segment)

    // ====================================================
    // 2. ��� ����
    // ====================================================

    // (1) Ŭ�� ���ֱ�
    clk_div u_clk_div (
        .clk(clk),
        .rst(rst),
        .o_tick(w_game_tick)
    );

    // (2) ���� Ÿ�̸�
    game_timer u_game_timer (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .cur_time(w_cur_time)
    );
    
    // (3) ��ư ��Ʈ�ѷ�
    button_ctrl u_btn_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_btn(i_btn),
        .o_start(w_start_btn), 
        .o_restart(w_restart_btn),
        .o_play(w_play_btn)
    );

    // (4) �Ǻ� FSM
    note_gen u_note_gen (
        .clk(clk),
        .rst(rst),
        .i_cur_time(w_cur_time),
        .o_note_t1(w_note_t1), 
        .o_note_t2(w_note_t2), 
        .o_game_end(w_game_end),
        .o_gen_pitch(w_gen_pitch)   // [����] ������ ����
    );
    
        // (7) LCD ��Ʈ�ѷ�
    lcd_ctrl u_lcd_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_note_t1(w_note_t1),
        .i_note_t2(w_note_t2),
        
        .o_lcd_rs(o_lcd_rs),
        .o_lcd_rw(o_lcd_rw),
        .o_lcd_e(o_lcd_e),
        .o_lcd_data(o_lcd_data),
        
        // ���� ��ȣ ����
        .o_hit_t1(w_hit_t1), 
        .o_hit_t2(w_hit_t2),
        
        .i_gen_pitch(w_gen_pitch),      // [����] ���� �޾Ƽ� ���
        .o_curr_pitch_t1(w_curr_pitch_t1), // [����] ��� �Ϸ�� ����
        .o_curr_pitch_t2(w_curr_pitch_t2)
    );
    
    // ���� ��Ʈ�ѷ�
    judgement_ctrl u_judge_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_btn_play(w_play_btn),
        .i_hit_t1(w_hit_t1),     // LCD ����
        .i_hit_t2(w_hit_t2),
        .i_curr_pitch_t1(w_curr_pitch_t1),
        .i_curr_pitch_t2(w_curr_pitch_t2),
        
        .o_judge(w_judge),
        .o_judge_hold(w_judge_hold),
        .o_play_en(w_play_en),   // -> Piezo �ѱ�
        .o_cnt_limit(w_cnt_limit) // -> Piezo ���ļ�
    );
    
    // ���� ���
    score_ctrl u_score_ctrl (
        .clk(clk),
        .rst(rst),
        .i_judge(w_judge),      // [�Է�] ���� ����� �޾Ƽ�
        .o_score(w_total_score) // [���] ���� ������ ����� ����
    );

    // Full Color LED
    full_color_led_ctrl u_led_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_game_over(w_game_end),
        .i_judge(w_judge_hold),      // [�Է�] ���� ����� �޾Ƽ� ���� ǥ��
        .o_fcl_r(o_fcl_r),
        .o_fcl_g(o_fcl_g),
        .o_fcl_b(o_fcl_b)
    );

    // ���� 7-Segment ��Ʈ�ѷ� (���� ���� 2,1,0 ǥ��)
    seven_segment_ctrl u_single_seg (
        .i_judge(w_judge_hold),      // ���� ��� �Է�
        .o_seg(o_single_seg)    // -> ���� ���׸�Ʈ ������ ���
    );

    // 8-Array Segment ��Ʈ�ѷ� (�ؽ�Ʈ + ���� ����)
    eight_array_seven_segment_ctrl u_array_seg (
        .clk(clk),
        .rst(rst),
        .i_judge(w_judge_hold),       // �ؽ�Ʈ ǥ�ÿ�
        .i_data(w_total_score),  // ���� ǥ�ÿ�
        .o_seg(o_array_seg),     // -> ��� ���׸�Ʈ ���� ��
        .o_com(o_array_com)      // -> ��� ���� ��
    );
    
    // (5) �ǿ��� ��Ʈ�ѷ�
    piezo_ctrl u_piezo_ctrl (
        .clk(clk), 
        .rst(rst), 
        .i_play_en(w_play_en),     // ���� ��⿡�� ���� ��ȣ�� �Ҹ� ��
        .i_cnt_limit(w_cnt_limit), // ���� ��⿡�� ���� ���ļ� ���
        .o_piezo(o_piezo)
    );

endmodule