module piezo_ctrl (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,
    input i_play_en,        // 1�� ���� �Ҹ� ��� (0�̸� ������)
    input [31:0] i_cnt_limit, // ���ļ� ������ ���� ī���� �� (�ܺο��� �־���)
    output reg o_piezo      // �ǿ��� ������ ������ ��ȣ
);

    reg [31:0] cnt;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            cnt <= 0;
            o_piezo <= 0;
        end else begin
            // �Ҹ� ��� �㰡(Enable)�� 1�� ���� ����
            if (i_play_en) begin
                // 6���� �ǽ� 2�� ���� ����
                // ī���Ͱ� ��ǥ��(���ֱ�)�� �����ϸ�
                if (cnt >= i_cnt_limit) begin
                    cnt <= 0;           // ī���� �ʱ�ȭ
                    o_piezo <= ~o_piezo; // ��ȣ ���� (0->1, 1->0)
                end else begin
                    cnt <= cnt + 1;     // ��� ��
                end
            end else begin
                // �Ҹ��� ����� �ϸ� �ʱ�ȭ
                cnt <= 0;
                o_piezo <= 0;
            end
        end
    end

endmodule