module intro_player (
    input clk,
    input rst,
    input i_tick,          // 1ms ƽ
    input i_enable,        // 1�� ���� �Ҹ� ��� (���� ���� ��)
    
    output reg o_play_en,      // �ǿ��� �ѱ�/����
    output reg [31:0] o_pitch  // �ǿ��� ���ļ� �� (Counter Limit)
);

    // ==========================================
    // "Sweet Child O' Mine" Riff Frequencies
    // ����: 50MHz / (Freq * 2)
    // ==========================================
    localparam D4  = 85132; // 293.66 Hz
    localparam D5  = 42565; // 587.33 Hz
    localparam A4  = 56818; // 440.00 Hz
    localparam G4  = 63775; // 392.00 Hz
    localparam G5  = 31888; // 783.99 Hz
    localparam Fs5  = 33784; // 739.99 Hz (F#5)

    // ���� ��Ʈ ���� (8�� �ݺ�)
    // Pattern: D4 -> D5 -> A4 -> G4 -> G5 -> A4 -> F#5 -> A4
    reg [31:0] riff_pitch [0:7];
    initial begin
        riff_pitch[0] = D4;
        riff_pitch[1] = D5;
        riff_pitch[2] = A4;
        riff_pitch[3] = G4;
        riff_pitch[4] = G5;
        riff_pitch[5] = A4;
        riff_pitch[6] = Fs5;
        riff_pitch[7] = A4;
    end

    // Ÿ�̹� ����
    parameter NOTE_DURATION = 200; // �� ���� 200ms (���� ���� ����)
    
    reg [31:0] time_cnt;
    reg [2:0]  note_idx; // 0~7

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            time_cnt <= 0;
            note_idx <= 0;
            o_play_en <= 0;
            o_pitch <= 0;
        end 
        else if (i_enable) begin
            // �Ҹ� �ѱ�
            o_play_en <= 1;
            o_pitch <= riff_pitch[note_idx];

            // Ÿ�̸� ����
            if (i_tick) begin
                if (time_cnt >= NOTE_DURATION - 1) begin
                    time_cnt <= 0;
                    note_idx <= note_idx + 1; // ���� ��Ʈ (�ڵ����� 0~7 �����÷ο�)
                end 
                else begin
                    time_cnt <= time_cnt + 1;
                end
            end
        end 
        else begin
            // ��Ȱ��ȭ �� �ʱ�ȭ
            o_play_en <= 0;
            o_pitch <= 0;
            time_cnt <= 0;
            note_idx <= 0;
        end
    end

endmodule