module sys_base (
    input clk,
    input rst
    // ... �ٸ� ����� ��Ʈ ...
);

    wire w_game_tick;      // �� ����� �̾��ִ� ����
    wire [31:0] w_cur_time; // ���� �ð��� ��� ����

    // ���ֱ� �ν��Ͻ� (Tick ����)
    clk_div u_clk_div (
        .clk(clk),
        .rst(rst),
        .o_tick(w_game_tick)
    );

    // Ÿ�̸� �ν��Ͻ� (�ð� ���)
    game_timer u_game_timer (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .cur_time(w_cur_time)
    );

    // ... ���� w_cur_time�� ����Ͽ� FSM ��� ���� ���� ���� ...

endmodule