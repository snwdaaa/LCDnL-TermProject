// Ŭ�� ���ֱ�
// �ٸ� ���鿡 1kHz Ŭ�� �Է�

module clk_div (
    input clk, // �ý��� Ŭ��
    input rst,
    output reg o_tick // ��� HIGH �Ǵ� tick ��ȣ
);

    // 100MHz -> 1kHz ��ȯ�� ���� ī���� ���Ѱ�
    // 100,000 - 1 = 99,999
    parameter CNT_MAX = 100000 - 1; 
    
    reg [31:0] cnt;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            cnt <= 0;
            o_tick <= 0;
        end else begin
            if (cnt >= CNT_MAX) begin
                cnt <= 0;
                o_tick <= 1; // 1ms �Ǹ� tick
            end else begin
                cnt <= cnt + 1;
                o_tick <= 0;
            end
        end
    end
endmodule