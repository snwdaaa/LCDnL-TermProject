`timescale 1ns / 1ps

module NOTE_GEN_TESTBENCH;

    // 1. �Է� ��ȣ (�츮�� ������ �͵�)
    reg clk;
    reg rst;
    reg [31:0] cur_time; // ��¥ ���� Ÿ�̸�

    // 2. ��� ��ȣ (������ �͵�)
    wire note_t1;    // ���� ��Ʈ ��ȣ
    wire note_t2;    // �Ʒ��� ��Ʈ ��ȣ
    wire game_end;   // ���� ���� ��ȣ

    // 3. ������ ���(DUT) ����
    note_gen u_note_gen (
        .clk(clk),
        .rst(rst),
        .i_cur_time(cur_time), // ���⿡ ��¥ �ð��� �ֽ��ϴ�
        .o_note_t1(note_t1),
        .o_note_t2(note_t2),
        .o_game_end(game_end)
    );

    // 4. Ŭ�� ���� (100MHz ����, �ֱ� 10ns)
    always #5 clk = ~clk;

    // 5. �׽�Ʈ �ó�����
    initial begin
        // �ʱ�ȭ
        clk = 0;
        rst = 1;
        cur_time = 0;

        // 1. ���� ����
        #20 rst = 0;
        
        // 2. �ð� ���� ����! (������ �ð��� �÷����ϴ�)
        $display("Start Simulation: Note Generation Test");

        // 0ms���� 8000ms���� 10ms ������ �ð��� ���� ������Ŵ
        // (���� ���Ӻ��� �ξ� ������ ������ �̴ϴ�)
        repeat (800) begin
            #10; // 10ns ��� (1Ŭ��)
            cur_time = cur_time + 10; // �ð��� 10ms�� �ǳʶ�
        end
        
        // 3. �ùķ��̼� ����
        #100;
        $display("Simulation Finish!");
        $finish;
    end

    // 6. ����͸� (�α� ���)
    // ��Ʈ ��ȣ�� 1�� �� ������ �ؽ�Ʈ�� �˷���
    always @(posedge clk) begin
        if (note_t1) 
            $display("[NOTE] Track 1 Fire! at Time: %d ms", cur_time);
        
        if (note_t2) 
            $display("[NOTE] Track 2 Fire! at Time: %d ms", cur_time);

        if (game_end)
            $display("[END] Game Over signal at Time: %d ms", cur_time);
    end

endmodule