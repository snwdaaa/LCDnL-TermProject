// ��Ʈ ������
// ���� ���� �ð��� ���� �Ǻ� ������ ���� ��ȣ ����

module note_gen (
    input clk,
    input rst,
    input [31:0] i_cur_time, // game_timer���� ���� ���� �ð� (ms)
    
    output reg o_note_t1,    // Track 1 (����) ��Ʈ ���� ��ȣ (1ƽ ���� 1)
    output reg o_note_t2,    // Track 2 (�Ʒ���) ��Ʈ ���� ��ȣ
    output reg [31:0] o_gen_pitch, // ������ ��Ʈ�� ���ļ� ��
    output reg o_game_end    // �뷡�� �������� �˸��� ��ȣ
);

    // Astronomia (Coffin Dance) Frequencies
    localparam F4  = 71586;  // �� (Main Base)
    localparam C5  = 47778;  // �� (High)
    localparam A4  = 56818;  // ��
    localparam G4  = 63775;  // ��
    localparam Bb4 = 53629;  // ��b
    localparam Ab4 = 60197;  // ��b (��#)
    localparam E4  = 75843;  // ��

    // ��Ʈ ���� ���� (16�� ���� * 8��Ʈ = 128��)
    parameter NOTE_COUNT = 200;
    integer i, j; // �ݺ��� ����
    
    // ���Ϻ� ���̽� ��Ʈ (ù 2�� ��) ����� �ӽ� ����
    reg [31:0] base_note;
    
    reg [31:0] note_time  [0:NOTE_COUNT-1];
    reg [1:0]  note_track [0:NOTE_COUNT-1];
    reg [31:0] note_pitch [0:NOTE_COUNT-1];
    
    // ���Ϻ� ���� �ð� ��� (�� ���ϴ� �� 1920ms)
    // idx: ���� ��Ʈ �ε��� (0 ~ 127)
    // time_offset: ���� ������ ���� �ð�
    integer idx;
    integer time_offset;

    initial begin
        // ==========================================
        // Megalovania (1�� ���� ����)
        // ==========================================
        
        // ��ü 4�� �ݺ� (1�� �� ������ 4���� ���� ����)
        for (i = 0; i < 4; i = i + 1) begin
            
            // 4���� ���� �ݺ� (D -> C -> B -> Bb)
            for (j = 0; j < 4; j = j + 1) begin
                
                idx = (i * 32) + (j * 8); 
                time_offset = 1000 + (i * 7680) + (j * 1920);

                // ���̽� ��Ʈ ���� (���ϸ��� �� 2�� ���� �ٸ�)
                if      (j == 0) base_note = D4;
                else if (j == 1) base_note = C4;
                else if (j == 2) base_note = B3;
                else             base_note = Bb3;

                // --- [Note 1] �� (Base) ---
                note_time [idx+0] = time_offset + 0;   note_track[idx+0] = 1; note_pitch[idx+0] = base_note;
                
                // --- [Note 2] �� (Base) ---
                note_time [idx+1] = time_offset + 120; note_track[idx+1] = 1; note_pitch[idx+1] = base_note; // ����!

                // --- [Note 3] �� (High D5) ---
                note_time [idx+2] = time_offset + 360; note_track[idx+2] = 2; note_pitch[idx+2] = D5; // ��Ÿ�� ����

                // --- [Note 4] �� (A4) ---
                note_time [idx+3] = time_offset + 600; note_track[idx+3] = 2; note_pitch[idx+3] = A4;
                
                // --- [Note 5] �� (Ab4) ---
                note_time [idx+4] = time_offset + 840; note_track[idx+4] = 1; note_pitch[idx+4] = Gs4;
                
                // --- [Note 6] �� (G4) ---
                note_time [idx+5] = time_offset + 1080; note_track[idx+5] = 2; note_pitch[idx+5] = G4;
                
                // --- [Note 7] �� (F4) ---
                note_time [idx+6] = time_offset + 1320; note_track[idx+6] = 1; note_pitch[idx+6] = F4;

                // --- [Note 8] ���� (D4 F4 G4) - ���⼭�� G4�� ������
                note_time [idx+7] = time_offset + 1560; note_track[idx+7] = 2; note_pitch[idx+7] = G4;
            end
        end
        
        // ������ ���� ó��
        // note_time[NOTE_COUNT] ó���� ���� (�ε��� ���� ��)
    end
    
    // ��Ʈ�� LCD ������ ���� �� �ɸ��� �ð� (�� 5�� ����)
    parameter END_DELAY = 5000;

    // ==========================================
    // ������ ���� (FSM)
    // ==========================================
    reg [31:0] note_idx; // ���� �� ��° ��Ʈ�� ��ٸ��� ������ (������)

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            note_idx <= 0;
            o_note_t1 <= 0;
            o_note_t2 <= 0;
            o_gen_pitch <= 0;
            o_game_end <= 0;
        end else begin
            o_note_t1 <= 0;
            o_note_t2 <= 0;

            // �뷡�� ���� �� �����ٸ�
            if (note_idx < NOTE_COUNT) begin
                // ���� �ð��� ��Ʈ�� �ð��� ���ų� ��������? (������ ��� ��� >= ���)
                if (i_cur_time >= note_time[note_idx]) begin
                    // ���� ���� ���
                    o_gen_pitch <= note_pitch[note_idx];
                    
                    // �ش� Ʈ���� ��ȣ �߻�
                    if (note_track[note_idx] == 1) 
                        o_note_t1 <= 1;
                    
                    if (note_track[note_idx] == 2) 
                        o_note_t2 <= 1;

                    // ���� ��Ʈ�� ������ �̵�
                    note_idx <= note_idx + 1;
                end
            end else begin
                // ��� ��Ʈ ���� ��, ������ ��Ʈ�� �������� ������ ������ ���
                // ex) ������ ��Ʈ �ð�(7700) + 5000ms = 12700ms�� �Ǿ�� ����
                if (i_cur_time >= note_time[NOTE_COUNT-1] + END_DELAY) begin
                    o_game_end <= 1;
                end
            end
        end
    end

endmodule