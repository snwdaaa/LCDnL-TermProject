module judgement_ctrl (
    input clk,
    input rst,
    input i_tick,           // 1ms ƽ (���� �ʱ�ȭ Ÿ�ֿ̹�)
    
    // �Է� ��ȣ
    input [1:0] i_btn_play, // [0]: Track 1 ��ư, [1]: Track 2 ��ư (ä�͸� ���ŵ�)

    // LCD ���� ��ȣ��
    input i_hit_t1,      // T1 Perfect Zone
    input i_pre_hit_t1,  // T1 Normal Zone
    input i_miss_t1,     // T1 Miss (������)
    
    input i_hit_t2,      // T2 Perfect Zone
    input i_pre_hit_t2,  // T2 Normal Zone
    input i_miss_t2,     // T2 Miss (������)
    
    input [31:0]  i_curr_pitch_t1,
    input [31:0] i_curr_pitch_t2,

    // ��� ��ȣ
    output reg [1:0] o_judge,      // ���� ��� (00:None, 11:Perfect ...)
    output reg [1:0] o_judge_hold, // [Hold]  ���÷��̿� (���� �������� ����) - NEW!
    output reg o_play_en,          // �ǿ��� �ѱ�
    output reg [31:0] o_cnt_limit, // �ǿ��� ���ļ� ��
    
    // ��Ʈ ���� ��û ��ȣ
    output reg o_clear_t1_perf,
    output reg o_clear_t1_norm,
    output reg o_clear_t2_perf,
    output reg o_clear_t2_norm
);

    // �Ҹ� ���� �ð��� ���� Ÿ�̸� (100ms)
    reg [31:0] sound_timer;
    parameter SOUND_DURATION = 100; // 100ms ���� ���

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_judge <= 0; o_judge_hold <= 0;
            o_play_en <= 0; o_cnt_limit <= 0;
            sound_timer <= 0;
            o_clear_t1_perf <= 0; o_clear_t1_norm <= 0;
            o_clear_t2_perf <= 0; o_clear_t2_norm <= 0;
        end else begin
            // Clear ��ȣ�� 1Ŭ���� �����ϰ� �ٷ� ���� �� (Pulse)
            o_clear_t1_perf <= 0; o_clear_t1_norm <= 0;
            o_clear_t2_perf <= 0; o_clear_t2_norm <= 0;

            // ====================================================
            // [Track 1 ����]
            // ====================================================
            if (i_btn_play[0]) begin
                // 1. Perfect (0�� ĭ)
                if (i_hit_t1) begin
                    o_judge <= 2'b11; o_judge_hold <= 2'b11; // Perfect
                    o_play_en <= 1; o_cnt_limit <= i_curr_pitch_t1;
                    sound_timer <= SOUND_DURATION;
                    o_clear_t1_perf <= 1; // ��Ʈ ���� ��û!
                end
                // 2. Normal (1�� ĭ) - Perfect�� �ƴ� ���� üũ
                else if (i_pre_hit_t1) begin
                    o_judge <= 2'b10; o_judge_hold <= 2'b10; // Normal
                    o_play_en <= 1; o_cnt_limit <= i_curr_pitch_t1; // (����� �ٻ�ġ ���)
                    sound_timer <= SOUND_DURATION;
                    o_clear_t1_norm <= 1; // ��Ʈ ���� ��û!
                end
            end
            
            // 3. Miss (��ư �� ������ ������)
            if (i_miss_t1) begin
                o_judge <= 2'b01; o_judge_hold <= 2'b01; // Miss
            end


            // ====================================================
            // [Track 2 ����] (���� ���� ����)
            // ====================================================
            if (i_btn_play[1]) begin
                if (i_hit_t2) begin
                    o_judge <= 2'b11; o_judge_hold <= 2'b11; 
                    o_play_en <= 1; o_cnt_limit <= i_curr_pitch_t2;
                    sound_timer <= SOUND_DURATION;
                    o_clear_t2_perf <= 1;
                end
                else if (i_pre_hit_t2) begin
                    o_judge <= 2'b10; o_judge_hold <= 2'b10; 
                    o_play_en <= 1; o_cnt_limit <= i_curr_pitch_t2;
                    sound_timer <= SOUND_DURATION;
                    o_clear_t2_norm <= 1;
                end
            end
            
            if (i_miss_t2) begin
                o_judge <= 2'b01; o_judge_hold <= 2'b01;
            end

            // ====================================================
            // ���� �ʱ�ȭ
            // ====================================================
            if (i_tick) begin
                o_judge <= 0; // ���� Pulse �ʱ�ȭ
                if (sound_timer > 0) sound_timer <= sound_timer - 1;
                else o_play_en <= 0;
            end
        end
    end

endmodule