module intro_player (
    input clk,
    input rst,
    input i_tick,          // 1ms ƽ (sys_base���� ������ Ÿ�̹� ��ȣ)
    input i_enable,        // 1�� ���� ���̷� �︲ (���� ���� �� or ���� ��)
    
    output reg o_play_en,      // �ǿ��� �ѱ�/����
    output reg [31:0] o_pitch  // �ǿ��� ���ļ� �� (Counter Limit)
);

    // ==========================================
    // ������ ���̷� ���ļ� ����
    // ����: 50MHz / (Freq * 2)
    // ==========================================
    // 400Hz (����) ~ 1000Hz (����) ���̸� �պ�
    localparam LOW_LIMIT  = 62500; // 400Hz
    localparam HIGH_LIMIT = 25000; // 1000Hz
    
    // �Ҹ� ��ȭ �ӵ� (���� Ŭ���� ������ ����)
    // 1ms���� �� ����ŭ ī���� ������ ���̰ų� �ø�
    localparam STEP = 25; 

    reg direction; // 0: ���� ������ (Limit ����), 1: ���� ������ (Limit ����)

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_pitch   <= LOW_LIMIT;
            direction <= 0;
            o_play_en <= 0;
        end 
        else if (i_enable) begin
            o_play_en <= 1; // �Ҹ� �ѱ�

            // 1ms���� ���ļ� ���� (�ε巯�� Sweep ȿ��)
            if (i_tick) begin
                if (direction == 0) begin 
                    // [��� ����] ��~~~~ (Limit ���� �ٿ��� ��������)
                    if (o_pitch > HIGH_LIMIT) 
                        o_pitch <= o_pitch - STEP;
                    else 
                        direction <= 1; // ���� ��ȯ (���� ��������)
                end 
                else begin 
                    // [�ϰ� ����] ��~~~~ (Limit ���� �÷��� ��������)
                    if (o_pitch < LOW_LIMIT) 
                        o_pitch <= o_pitch + STEP;
                    else 
                        direction <= 0; // ���� ��ȯ (���� �ö���)
                end
            end
        end 
        else begin
            // ��Ȱ��ȭ �� (���� ���� ��) �Ҹ� ���� �ʱ�ȭ
            o_play_en <= 0;
            o_pitch   <= LOW_LIMIT; 
            direction <= 0;
        end
    end

endmodule