module u_game_8a_7_segment (
    input clk,
    input rst,
    input [1:0] i_judge,    // 00:IDLE, 01:MISS, 10:NORMAL, 11:PERFECT
    output reg [7:0] o_seg, // Segment Pattern (a~g, dp)
    output reg [7:0] o_com  // Digit Selection (Active Low)
);

    // [1] ���� ���� ���� (Active Low: 0�� �� ����)
    // a=MSB(7), dp=LSB(0) �Ǵ� a=0, dp=7 �� ���帶�� �ٸ�. 
    // ���⼭�� �Ϲ����� [7:0] = {dp, g, f, e, d, c, b, a} ���� Ȥ�� ���� �޴��� ����.
    // �� HBE-Combo II ���� Ư���� ���� a(bit0)~g(bit6), dp(bit7)�� �����ϰ�, 0=ON���� �����մϴ�.
    // ��Ʈ ������ �ٸ��� .xdc ���Ͽ��� ������ �ٲٰų� ���⼭ ���� �������� �˴ϴ�.
    
    localparam CH_BLK = 8'b1111_1111; // ���� (Blank)
    localparam CH_P   = 8'b0000_1100; // P
    localparam CH_E   = 8'b0000_0110; // E
    localparam CH_R   = 8'b1010_1111; // r (�ҹ��� ���)
    localparam CH_F   = 8'b0000_1110; // F
    localparam CH_C   = 8'b0100_0110; // C
    localparam CH_T   = 8'b0000_0111; // t
    localparam CH_N   = 8'b1010_1011; // n
    localparam CH_O   = 8'b1010_0011; // o
    localparam CH_M   = 8'b1010_1010; // n �ΰ� ��ģ ��� (M�� ǥ���� ����� �ٻ�ġ ���)
    localparam CH_I   = 8'b1111_1001; // I (1�� ����)
    localparam CH_S   = 8'b0001_0010; // S (5�� ����)
    localparam CH_A   = 8'b0000_1000; // A
    localparam CH_L   = 8'b1000_0111; // L

    // [2] ��ĳ�� Ÿ�̸� (Scanning Timer)
    // 8�� �ڸ��� ������ ��ȯ�ϱ� ���� ī����
    reg [16:0] scan_cnt;
    always @(posedge clk or posedge rst) begin
        if (rst) scan_cnt <= 0;
        else scan_cnt <= scan_cnt + 1;
    end
    
    // ���� 3��Ʈ�� ����Ͽ� 0~7�� �ڸ��� ��ȯ (2^3 = 8��)
    wire [2:0] scan_idx = scan_cnt[16:14];

    // [3] �ڸ��� ���� �� ���� ��� ����
    // scan_idx(���� ���� �ڸ�)�� i_judge(���� ����)�� ���� ����� ���� ����
    // �ڸ� ��ġ: scan_idx 7(����/MSB) -> 0(������/LSB)
    always @(*) begin
        // 1. Common �� ���� (Active Low) - ���� scan_idx�� �ش��ϴ� �ڸ��� 0����
        o_com = ~(8'b0000_0001 << scan_idx); 

        // 2. Segment ������ ����
        case (i_judge)
            // -----------------------------------------------------
            // Case 1: PERFECT ( "P E r F E C t _" )
            // -----------------------------------------------------
            2'b11: begin 
                case (scan_idx)
                    3'd7: o_seg = CH_P;   // [7] P
                    3'd6: o_seg = CH_E;   // [6] E
                    3'd5: o_seg = CH_R;   // [5] r
                    3'd4: o_seg = CH_F;   // [4] F
                    3'd3: o_seg = CH_E;   // [3] E
                    3'd2: o_seg = CH_C;   // [2] C
                    3'd1: o_seg = CH_T;   // [1] t
                    default: o_seg = CH_BLK; // ������ ����
                endcase
            end

            // -----------------------------------------------------
            // Case 2: NORMAL ( "n o r n A L _ _" )
            // -----------------------------------------------------
            2'b10: begin
                case (scan_idx)
                    3'd7: o_seg = CH_N;   // [7] n
                    3'd6: o_seg = CH_O;   // [6] o
                    3'd5: o_seg = CH_R;   // [5] r
                    3'd4: o_seg = CH_N;   // [4] n
                    3'd3: o_seg = CH_A;   // [3] A
                    3'd2: o_seg = CH_L;   // [2] L
                    default: o_seg = CH_BLK; // ������ ����
                endcase
            end

            // -----------------------------------------------------
            // Case 3: MISS ( "_ _ n I S S _ _" ) - �߾� ���� ����
            // -----------------------------------------------------
            2'b01: begin
                case (scan_idx)
                    3'd5: o_seg = CH_N;   // [5] M (n ��� ���)
                    3'd4: o_seg = CH_I;   // [4] I
                    3'd3: o_seg = CH_S;   // [3] S
                    3'd2: o_seg = CH_S;   // [2] S
                    default: o_seg = CH_BLK; // ������ ����
                endcase
            end

            // -----------------------------------------------------
            // Case 0: IDLE ( "_ _ _ _ _ _ _ _" )
            // -----------------------------------------------------
            default: o_seg = CH_BLK; // �ƹ��͵� ǥ�� �� ��
        endcase
    end

endmodule