module sys_base (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,              // ����
    
    // �ǿ��� ���� ��� (������ ���� �ǵ��)
    output o_piezo,
    
    // LCD ���� ��
    output o_lcd_rs,
    output o_lcd_rw,
    output o_lcd_e,
    output [7:0] o_lcd_data,
    
    // ��ư �Է�
    input [3:0] i_btn       // ��ư �Է� 4��
);

    // ====================================================
    // 1. ���� ��ȣ ����
    // ====================================================
    wire w_game_tick;       // 1ms ƽ
    wire [31:0] w_cur_time; // ���� ���� �ð�
    
    // ��Ʈ ��ȣ
    wire w_note_t1;         // ���� ��Ʈ
    wire w_note_t2;         // �Ʒ��� ��Ʈ
    wire w_game_end;
    
    // ��ư ��ȣ (ä�͸� ���ŵ�)
    wire w_start_btn;
    wire w_restart_btn;
    wire [1:0] w_play_btn;  // [1]: Down(Track2), [0]: Up(Track1)
    
    // �ǿ��� ���� ��ȣ (Judgement -> Piezo)
    wire w_play_en;         // �Ҹ� ��� Enable
    wire [31:0] w_cnt_limit;// ����� ���ļ� ��
    
    // ���� ��� ��ȣ (���� ��� �� ��, ���� Ȯ���)
    wire [1:0] w_judge;     
    
    // LCD ������ ���� ��ȣ
    wire w_hit_t1, w_hit_t2;

    // ====================================================
    // 2. ��� ����
    // ====================================================

    // (1) Ŭ�� ���ֱ�
    clk_div u_clk_div (
        .clk(clk),
        .rst(rst),
        .o_tick(w_game_tick)
    );

    // (2) ���� Ÿ�̸�
    game_timer u_game_timer (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .cur_time(w_cur_time)
    );
    
    // (3) ��ư ��Ʈ�ѷ�
    button_ctrl u_btn_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_btn(i_btn),
        .o_start(w_start_btn), 
        .o_restart(w_restart_btn),
        .o_play(w_play_btn)
    );

    // (4) �Ǻ� FSM
    note_gen u_note_gen (
        .clk(clk),
        .rst(rst),
        .i_cur_time(w_cur_time),
        .o_note_t1(w_note_t1), 
        .o_note_t2(w_note_t2), 
        .o_game_end(w_game_end)
    );
    
    // (5) �ǿ��� ��Ʈ�ѷ�
    piezo_ctrl u_piezo_ctrl (
        .clk(clk), 
        .rst(rst), 
        .i_play_en(w_play_en),     // ���� ��⿡�� ���� ��ȣ�� �Ҹ� ��
        .i_cnt_limit(w_cnt_limit), // ���� ��⿡�� ���� ���ļ� ���
        .o_piezo(o_piezo)
    );
    
    // (6) ���� ��Ʈ�ѷ�
    judgement_ctrl u_judge_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_btn_play(w_play_btn),
        .i_hit_t1(w_hit_t1),     // LCD ����
        .i_hit_t2(w_hit_t2),
        
        .o_judge(w_judge),
        .o_play_en(w_play_en),   // -> Piezo �ѱ�
        .o_cnt_limit(w_cnt_limit) // -> Piezo ���ļ�
    );

    // (7) LCD ��Ʈ�ѷ�
    lcd_ctrl u_lcd_ctrl (
        .clk(clk),
        .rst(rst),
        .i_tick(w_game_tick),
        .i_note_t1(w_note_t1),
        .i_note_t2(w_note_t2),
        
        .o_lcd_rs(o_lcd_rs),
        .o_lcd_rw(o_lcd_rw),
        .o_lcd_e(o_lcd_e),
        .o_lcd_data(o_lcd_data),
        
        // ���� ��ȣ ����
        .o_hit_t1(w_hit_t1), 
        .o_hit_t2(w_hit_t2)
    );

endmodule