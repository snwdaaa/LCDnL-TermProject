module score_ctrl (
    input clk,
    input rst,
    input [1:0] i_judge,     // ���� ��� (11:Perfect, 10:Normal, 01:Miss)
    output reg [15:0] o_score // ������ �� ����
);

    reg [1:0] judge_prev;    // ���� ���ؼǿ� ���� ���� ����

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_score <= 0;
            judge_prev <= 0;
        end else begin
            judge_prev <= i_judge;

            // [�ٽ�] ���� ��ȣ�� ���ϴ� ����(Rising Edge)���� ���� �ջ�
            // 00(Idle)�� �ƴϰ�, ���� ���¿� �ٸ� �� ����
            if (i_judge != 0 && i_judge != judge_prev) begin
                case (i_judge)
                    2'b11: o_score <= o_score + 2; // Perfect: +2��
                    2'b10: o_score <= o_score + 1; // Normal: +1��
                    2'b01: o_score <= o_score + 0; // Miss: +0��
                    default: ;
                endcase
            end
        end
    end
endmodule