module lcd_ctrl (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,              // ����
    input i_tick,           // 1ms ƽ (��ũ�� �ӵ� ������)
    
    // ��Ʈ ���� ��ȣ (from note_gen)
    // 1Ŭ�� ���ȸ� '��¦'�ϹǷ� ��ġ�� �ʰ� ��ƾ� �մϴ�.
    input i_note_t1,        // ���� (Track 1) ��Ʈ
    input i_note_t2,        // �Ʒ��� (Track 2) ��Ʈ
    
    input [31:0] i_gen_pitch, // note_gen���� ���� ����
    
    // LCD �ϵ���� �� (���� �ɿ� ����)
    output reg o_lcd_rs,    // 0:���, 1:������
    output reg o_lcd_rw,    // 0:����, 1:�б� (�׻� 0)
    output reg o_lcd_e,     // Enable �޽�
    output reg [7:0] o_lcd_data, // ������ ����
    
    // ������(�� ����) ���� �˸� ��ȣ
    output o_hit_t1, // Track 1 �������� ��Ʈ ����!
    output o_hit_t2,  // Track 2 �������� ��Ʈ ����!
    
    // ���� �������� �ִ� ��Ʈ�� ���� ��
    output reg [31:0] o_curr_pitch_t1, 
    output reg [31:0] o_curr_pitch_t2
);

    // ====================================================
    // [Part 1] ��Ʈ ��ũ�Ѹ� ���� (Buffer & Scroll)
    // ====================================================
    
    // 1. ȭ�� ���� (16ĭ x 2��)
    reg [7:0] line1 [0:15]; // ����
    reg [7:0] line2 [0:15]; // �Ʒ���
    
    // ���� ���� (ȭ��� �Ȱ��� �̵��ϴ� ������ ������ ����)
    reg [31:0] pitch_buf_t1 [0:15];
    reg [31:0] pitch_buf_t2 [0:15];

    // 2. ��Ʈ ĸó (Note Capture)
    // note_gen���� ������ ��ȣ�� ���� ª���Ƿ�(1Ŭ��), 
    // ���� ��ũ���� �Ͼ ������ ����ص־� �մϴ�.
    reg r_catch_t1, r_catch_t2;
    
    // ĸó�� ��������
    reg [31:0] r_catch_pitch;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            r_catch_t1 <= 0; r_catch_t2 <= 0;
            r_catch_pitch <= 0;
        end else begin
            if (i_note_t1) begin
                    r_catch_t1 <= 1;
                    r_catch_pitch <= i_gen_pitch; // ���赵 ���� ĸó!
            end else if (scroll_en) r_catch_t1 <= 0; // ��ũ�� �� �ʱ�ȭ
            
            if (i_note_t2) begin
                r_catch_t2 <= 1;
                r_catch_pitch <= i_gen_pitch;
            end else if (scroll_en) r_catch_t2 <= 0;
        end
    end

    // 3. ��ũ�� Ÿ�̸� (Scroll Timer)
    // 300ms���� �� ĭ�� �̵� (�ӵ� ���� ����)
    parameter SCROLL_SPEED = 300; 
    reg [31:0] scroll_cnt;
    wire scroll_en;

    always @(posedge clk or posedge rst) begin
        if (rst) scroll_cnt <= 0;
        else if (i_tick) begin
            if (scroll_cnt >= SCROLL_SPEED - 1) scroll_cnt <= 0;
            else scroll_cnt <= scroll_cnt + 1;
        end
    end
    assign scroll_en = (i_tick && (scroll_cnt == 0));

    // 4. ���� ������Ʈ (Shift Logic)
    integer i;
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            // �ʱ�ȭ: ����(" ")���� ä�� (ASCII 0x20)
            for (i=0; i<16; i=i+1) begin
                line1[i] <= 8'h20;
                line2[i] <= 8'h20;
                
                // ���赵 �Ȱ��� �ʱ�ȭ
                pitch_buf_t1[i] <= 0;
                pitch_buf_t2[i] <= 0;
            end
        end else if (scroll_en) begin
            // [�������� �̵�]
            for (i=0; i<15; i=i+1) begin
                line1[i] <= line1[i+1];
                line2[i] <= line2[i+1];
                
                // ���赵 �Ȱ��� �̵�
                pitch_buf_t1[i] <= pitch_buf_t1[i+1];
                pitch_buf_t2[i] <= pitch_buf_t2[i+1];
            end
            
            // [������ �� ä���]
            // ��Ҵ� ��Ʈ�� ������ 'O' (0x4F), ������ ���� ' ' (0x20)
            line1[15] <= (r_catch_t1) ? 8'h4F : 8'h20;
            line2[15] <= (r_catch_t2) ? 8'h4F : 8'h20;
            pitch_buf_t1[15] <= (r_catch_t1) ? r_catch_pitch : 0;
            pitch_buf_t2[15] <= (r_catch_t2) ? r_catch_pitch : 0;
        end
    end
    
    // [Part 3] ������ ���� ��� (�� �Ʒ��� �߰��ϼ���!)
    // �� ����(0��) ĭ ���� ���� 'O'(0x4F)�̸� 1�� ����մϴ�.
    assign o_hit_t1 = (line1[0] == 8'h4F);
    assign o_hit_t2 = (line2[0] == 8'h4F);
    
    // �� ����(0��) ĭ�� ������ �������ϴ�.
    always @(*) begin
        o_curr_pitch_t1 = pitch_buf_t1[0];
        o_curr_pitch_t2 = pitch_buf_t2[0];
    end

    // ====================================================
    // [Part 2] LCD ����̹� (Hardware Control FSM)
    // ====================================================
    
    // ���� ����
    localparam S_INIT       = 0; // �ʱ�ȭ ���
    localparam S_CMD_PRE    = 1; // ��� ���� �غ�
    localparam S_CMD_SEND   = 2; // ��� ���� (E=1)
    localparam S_CMD_HOLD   = 3; // ��� �Ϸ� ���
    localparam S_DATA_PRE   = 4; // ������ ���� �غ�
    localparam S_DATA_SEND  = 5; // ������ ���� (E=1)
    localparam S_DATA_HOLD  = 6; // ������ �Ϸ� ���
    
    reg [3:0] state;
    reg [4:0] init_step;     // �ʱ�ȭ �ܰ�
    reg [4:0] char_idx;      // ���� ���� �ִ� ���� ��ġ (0~31)
    
    reg [31:0] delay_cnt;    // Ÿ�̹� ���߱� ���� ī����
    
    // 50MHz Ŭ�� ���� ������ ���
    // 2ms = 100,000 Ŭ�� (Clear �� �� ���)
    // 50us = 2,500 Ŭ�� (�Ϲ� ���)
    parameter DLY_2MS = 100000;
    parameter DLY_50US = 2500;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= S_INIT;
            init_step <= 0;
            char_idx <= 0;
            delay_cnt <= 0;
            o_lcd_e <= 0;
            o_lcd_rs <= 0;
            o_lcd_rw <= 0;
            o_lcd_data <= 0;
        end else begin
            case (state)
                // ------------------------------------------------
                // 1. �ʱ�ȭ (Initialization Sequence)
                // ------------------------------------------------
                S_INIT: begin
                    delay_cnt <= delay_cnt + 1;
                    // ���� �Ѱ� ����� ��ٸ� (�� 15ms �̻� -> �˳��� 20ms)
                    if (delay_cnt > DLY_2MS * 10) begin 
                        delay_cnt <= 0;
                        state <= S_CMD_PRE;
                    end
                end

                // ------------------------------------------------
                // 2. ��� ������ (Command Send)
                // ------------------------------------------------
                S_CMD_PRE: begin
                    o_lcd_rs <= 0; // ��� ���
                    o_lcd_rw <= 0; // ����
                    o_lcd_e  <= 0;
                    
                    // �ʱ�ȭ �ܰ躰 ��ɾ� ����
                    case (init_step)
                        0: o_lcd_data <= 8'h38; // Function Set (8bit, 2line)
                        1: o_lcd_data <= 8'h0C; // Display ON, Cursor OFF
                        2: o_lcd_data <= 8'h06; // Entry Mode (Auto Inc)
                        3: o_lcd_data <= 8'h01; // Clear Display
                        4: o_lcd_data <= 8'h80; // Line 1 ���� �ּ� (0x80)
                        5: o_lcd_data <= 8'hC0; // Line 2 ���� �ּ� (0xC0)
                        default: o_lcd_data <= 8'h80; // (Refresh Loop ����)
                    endcase
                    state <= S_CMD_SEND;
                end

                S_CMD_SEND: begin
                    o_lcd_e <= 1; // Enable Pulse High
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > 50) begin // ������ �޽� �� ����
                        delay_cnt <= 0;
                        state <= S_CMD_HOLD;
                    end
                end
                
                S_CMD_HOLD: begin
                    o_lcd_e <= 0; // Enable Pulse Low
                    delay_cnt <= delay_cnt + 1;
                    
                    // Clear ���(step 3)�� ���� �ɸ� (2ms), �������� ���� (50us)
                    if ((init_step == 3 && delay_cnt > DLY_2MS) || 
                        (init_step != 3 && delay_cnt > DLY_50US)) begin
                        
                        delay_cnt <= 0;
                        
                        // �ʱ�ȭ ���̸� ���� �ܰ��
                        if (init_step < 4) begin
                            init_step <= init_step + 1;
                            state <= S_CMD_PRE;
                        end 
                        // �ʱ�ȭ �������� ������ ���� ����
                        else begin
                            // ȭ�� ���� ����: Line 1 �ּ� ����(4) -> Line 1 ������ ����
                            // -> Line 2 �ּ� ����(5) -> Line 2 ������ ����
                            if (init_step == 4) begin
                                char_idx <= 0;      // 0~15�� ���� �� �غ�
                                state <= S_DATA_PRE; 
                            end else if (init_step == 5) begin
                                char_idx <= 16;     // 16~31�� ���� �� �غ�
                                state <= S_DATA_PRE;
                            end
                        end
                    end
                end

                // ------------------------------------------------
                // 3. ������ ������ (Data Send - ȭ�� �׸���)
                // ------------------------------------------------
                S_DATA_PRE: begin
                    o_lcd_rs <= 1; // ������ ���
                    o_lcd_rw <= 0;
                    o_lcd_e  <= 0;
                    
                    // ���� char_idx�� �´� ���� ���� ��������
                    if (char_idx < 16) 
                        o_lcd_data <= line1[char_idx];      // ����
                    else 
                        o_lcd_data <= line2[char_idx - 16]; // �Ʒ���
                        
                    state <= S_DATA_SEND;
                end

                S_DATA_SEND: begin
                    o_lcd_e <= 1;
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > 50) begin
                        delay_cnt <= 0;
                        state <= S_DATA_HOLD;
                    end
                end

                S_DATA_HOLD: begin
                    o_lcd_e <= 0;
                    delay_cnt <= delay_cnt + 1;
                    if (delay_cnt > DLY_50US) begin // 50us ���
                        delay_cnt <= 0;
                        
                        // ���� ���ڷ� �̵�
                        if (char_idx == 15) begin
                            // ���� �� ������ -> �Ʒ��� �ּ� �����Ϸ� ����
                            init_step <= 5; 
                            state <= S_CMD_PRE;
                        end else if (char_idx == 31) begin
                            // �Ʒ��� �� ������ -> �ٽ� ���� �ּ� �����Ϸ� ���� (���� ����)
                            init_step <= 4; 
                            state <= S_CMD_PRE;
                        end else begin
                            // ���� �� ���� ����
                            char_idx <= char_idx + 1;
                            state <= S_DATA_PRE;
                        end
                    end
                end
            endcase
        end
    end

endmodule