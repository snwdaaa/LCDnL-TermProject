`timescale 1ns / 1ps

module CLK_TESTBENCH;

    // 1. �Է� ��ȣ ���� (reg)
    reg clk;
    reg rst;

    // 2. ������ ���(DUT) �ν��Ͻ� ����
    sys_base u_sys_base (
        .clk(clk),
        .rst(rst)
    );

    // 3. 50MHz Ŭ�� ���� (�ֱ� 20ns)
    // 10ns���� ���� �������� �ֱ�� 20ns�� �˴ϴ�.
    always #10 clk = ~clk;

    // 4. �׽�Ʈ �ó�����
    initial begin
        // �ʱ�ȭ
        clk = 0;
        rst = 1; // ���� �� ������

        // �ùķ��̼� ���� �޽���
        $display("Simulation Start!");

        // 100ns �� ���� ���� (���� ����)
        #100;
        rst = 0;
        $display("Reset released. Game Timer should start counting...");

        // ����� �ð� ���� �ùķ��̼� ����
        // ����: CNT_MAX�� ������ �ʾҴٸ� 1ms�� ���� ���� �ſ� ���� ������ �մϴ�.
        // ���⼭�� ���÷� 5000ns�� �����ϴ�.
        #5000;

        $display("Simulation Finish!");
        $finish;
    end
    
    // 5. ����͸� (�ɼ�)
    // �ùķ��̼� �α�â�� ���� �ؽ�Ʈ�� ���� �ʹٸ� �Ʒ� ���� Ȱ��
    // u_sys_base ������ u_game_timer ����� cur_time ���� ���ĺ��ϴ�.
    always @(posedge clk) begin
        // ���� ���� ������ �α� ��� (Hierarchical Reference ���)
        if (u_sys_base.w_game_tick) begin
            $display("Time: %d ms", u_sys_base.w_cur_time);
        end
    end

endmodule