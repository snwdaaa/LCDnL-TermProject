module led_ctrl (
    input clk,              // �ý��� Ŭ�� (50MHz)
    input rst,              // ����
    input i_tick,           // 1ms ƽ (�ӵ� ������)
    input i_game_start,     // ���� ���� ��ȣ (1�� ���� ������)
    input i_game_over,      // (����) ���� ���� �� �����̰� �� ���� ����
    
    output reg [7:0] o_led  // 8�� LED ���
);

    // ==========================================
    // ����: �ӵ� ����
    // ==========================================
    parameter MOVE_SPEED = 100; // 100ms���� �� ĭ �̵� (�������� ����)
    
    reg [31:0] move_cnt;    // �ð� ī����
    reg [2:0]  led_idx;     // ���� ���� LED ��ġ (0~7)
    reg        dir;         // �̵� ���� (0: ����->������, 1: ������->����)

    // ==========================================
    // ���� ����
    // ==========================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_led <= 8'b0000_0000;
            move_cnt <= 0;
            led_idx <= 0;
            dir <= 0;
        end 
        else if (i_game_start && !i_game_over) begin
            // 1. Ÿ�̸� ���� (MOVE_SPEED ���� Ʈ����)
            if (i_tick) begin
                if (move_cnt >= MOVE_SPEED - 1) begin
                    move_cnt <= 0;
                    
                    // 2. LED ��ġ �̵� �� ���� ��ȯ
                    if (dir == 0) begin 
                        // [������] 0 -> 7
                        if (led_idx == 7) begin
                            dir <= 1;       // ���� ������ ���� �ݴ��
                            led_idx <= 6;
                        end else begin
                            led_idx <= led_idx + 1;
                        end
                    end 
                    else begin 
                        // [������] 7 -> 0
                        if (led_idx == 0) begin
                            dir <= 0;       // ���� ������ ���� �ݴ��
                            led_idx <= 1;
                        end else begin
                            led_idx <= led_idx - 1;
                        end
                    end
                end 
                else begin
                    move_cnt <= move_cnt + 1;
                end
            end
            
            // 3. ���� ��ġ�� LED �ѱ� (Decoder)
            o_led <= (8'b1 << led_idx);
            
        end 
        else begin
            // ���� ���� �ƴ� ���� ��� ���ų�, Ư�� ���� ����
            o_led <= 8'b0000_0000;
            move_cnt <= 0;
            led_idx <= 0;
        end
    end

endmodule