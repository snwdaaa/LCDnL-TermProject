module u_game_button (
    input clk,              // �ý��� Ŭ��
    input rst,              // ����
    input i_tick,           // 1ms ƽ (��ٿ�� �ð� ������)
    input [3:0] i_btn,      // ���� ������ ��ư �Է� (4��)
    
    // ������ ��� ��ȣ (���Һ� �и�)
    output o_start,         // ���� ���� (One-shot)
    output o_restart,       // ���� ����� (One-shot)
    output [1:0] o_play     // �÷��� ��ư 2�� (One-shot)
);

    // [1] ��ư ���� ���� (����ϱ� ���ϰ� �ε��� ����)
    // ������ ��ư ������ ���� ������ ������ �� �ֽ��ϴ�.
    localparam IDX_START   = 0;
    localparam IDX_RESTART = 1;
    localparam IDX_PLAY_L  = 2;
    localparam IDX_PLAY_R  = 3;

    // [2] ���� �������� ����
    reg [3:0] btn_stable;   // ��ٿ���� �Ϸ�� �������� ����
    reg [3:0] btn_prev;     // ���� ������ ���� ���� ���� ����
    
    // �� ��ư���� ä�͸��� �Ÿ��� ���� ī���� (4��)
    reg [4:0] debounce_cnt [0:3]; 
    parameter DEBOUNCE_TIME = 20; // 20ms ���� ��ȣ�� �����Ǿ�� ����

    integer i;

    // [3] ��ٿ�� ���� (Debouncing)
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            btn_stable <= 4'b0000;
            for (i=0; i<4; i=i+1) debounce_cnt[i] <= 0;
        end else if (i_tick) begin
            for (i=0; i<4; i=i+1) begin
                // �Է�(i_btn)�� ���� ������ ����(btn_stable)�� �ٸ��� ī��Ʈ ����
                if (i_btn[i] != btn_stable[i]) begin
                    if (debounce_cnt[i] >= DEBOUNCE_TIME - 1) begin
                        btn_stable[i] <= i_btn[i]; // 20ms ��� �� ���� ������Ʈ
                        debounce_cnt[i] <= 0;
                    end else begin
                        debounce_cnt[i] <= debounce_cnt[i] + 1;
                    end
                end else begin
                    debounce_cnt[i] <= 0; // ������ٸ� ī���� �ʱ�ȭ
                end
            end
        end
    end

    // [4] ���� ���� ���� (Edge Detection)
    // ��ư�� 0 -> 1�� ���ϴ� ����(Rising Edge)�� 1�� ���
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            btn_prev <= 4'b0000;
        end else begin
            btn_prev <= btn_stable;
        end
    end

    // ����� 1�̰�, ������ 0�̾��� ���� (Rising Edge)
    wire [3:0] btn_rise = btn_stable & ~btn_prev;

    // [5] ��� �Ҵ� (���� �й�)
    assign o_start   = btn_rise[IDX_START];
    assign o_restart = btn_rise[IDX_RESTART];
    assign o_play    = {btn_rise[IDX_PLAY_R], btn_rise[IDX_PLAY_L]};

endmodule