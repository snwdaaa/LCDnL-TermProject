module u_game_led (
    input clk,              // �ý��� Ŭ�� (100MHz or 50MHz)
    input rst,              // ���� ��ȣ
    input i_tick,           // 1ms ƽ (clk_div ��⿡�� �޾ƿ�)
    input i_spawn_note,     // ��Ʈ ���� ��ȣ (1 = ��Ʈ ����, �Ǻ� or ��ư���� �Է�)
    output reg [7:0] o_led, // LED ��� (�̰� ���� LED �ɿ� ����)
    output o_is_target      // [�߿�] Ÿ��(LED8) ���� �˸� ��ȣ (���߿� ���� ��⿡ ����)
);

    // [1] �ӵ� ���� �Ķ���� (���̵� ����)
    // 200 = 200ms���� �� ĭ �̵�. ���ڸ� ���̸� �������ϴ�.
    parameter NOTE_SPEED = 200; 

    reg [31:0] speed_cnt;
    wire move_en; // �̵� �㰡 ��ȣ

    // [2] �̵� Ÿ�̹� ���� ���� (Timer)
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            speed_cnt <= 0;
        end else if (i_tick) begin
            // NOTE_SPEED ��ŭ 1ms ƽ�� ���ϴ�.
            if (speed_cnt >= NOTE_SPEED - 1) begin
                speed_cnt <= 0;
            end else begin
                speed_cnt <= speed_cnt + 1;
            end
        end
    end

    // ī���Ͱ� 0�� �Ǵ� �������� 1������ High�� �˴ϴ�.
    assign move_en = (i_tick && (speed_cnt == 0));

    // [3] ����Ʈ �������� ���� (�ٽ�: ������ �̵�)
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_led <= 8'b00000000; // �ʱ�ȭ: ��� �� ����
        end else if (move_en) begin
            // [�̵� ����: Left -> Right]
            // o_led ���� �������� Shift (<< 1) �Ͽ� �����͸� ���� ��Ʈ�� �Ӵϴ�.
            // �� �ڸ��� �� 0�� ��Ʈ(LSB) �ڸ��� i_spawn_note ���� ä�� �ֽ��ϴ�.
            // ��: 00000000 -> 00000001 -> 00000010 -> ... -> 10000000
            o_led <= (o_led << 1) | i_spawn_note;
        end
    end

    // [4] Ÿ�� ���� Ȯ��
    // ���� ������(LED8)�� 7�� ��Ʈ�� ���� ���Դ��� Ȯ��
    assign o_is_target = o_led[7]; 

endmodule