// ���ֱ⿡�� ���� tick ��ȣ �޾Ƽ�
// ���� ���� �� �� �� ms �������� ���� �ð� ��

module game_timer (
    input clk, // �ý��� Ŭ��
    input rst,
    input i_tick, // ���ֱ⿡�� ���� 1ms ƽ ��ȣ
    output reg [31:0] cur_time // ���� ���� �ð� (ms ����)
);

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            cur_time <= 0;
        end else begin
            if (i_tick) begin
                cur_time <= cur_time + 1; // 1ms ƽ�� ���� ���� �ð� ����
            end
        end
    end
endmodule