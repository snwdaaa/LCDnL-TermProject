module judgement_ctrl (
    input clk,
    input rst,
    input i_tick,           // 1ms ƽ (���� �ʱ�ȭ Ÿ�ֿ̹�)
    
    // �Է� ��ȣ
    input [1:0] i_btn_play, // [0]: Track 1 ��ư, [1]: Track 2 ��ư (ä�͸� ���ŵ�)
    input i_hit_t1,         // Track 1 ������ ���� (LCD���� ��)
    input i_hit_t2,         // Track 2 ������ ���� (LCD���� ��)
    
    input [31:0]  i_curr_pitch_t1,
    input [31:0] i_curr_pitch_t2,

    // ��� ��ȣ
    output reg [1:0] o_judge,      // ���� ��� (00:None, 11:Perfect ...)
    output reg o_play_en,          // �ǿ��� �ѱ�
    output reg [31:0] o_cnt_limit // �ǿ��� ���ļ� ��
);

    // �Ҹ� ���� �ð��� ���� Ÿ�̸� (100ms)
    reg [31:0] sound_timer;
    parameter SOUND_DURATION = 100; // 100ms ���� ���

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            o_judge <= 0;
            o_play_en <= 0;
            o_cnt_limit <= 0;
            sound_timer <= 0;
        end else begin
            // ====================================================
            // 1. ���� ���� (Priority: Track 1 -> Track 2)
            // ====================================================
            
            // [Track 1 ����?] LCD�� ��Ʈ �ְ�(i_hit_t1) & ��ư ������ ��(i_btn_play[0])
            if (i_hit_t1 && i_btn_play[0]) begin
                o_judge <= 2'b11;        // Perfect!
                o_play_en <= 1;          // �Ҹ� ON
                o_cnt_limit <= i_curr_pitch_t1;  // LCD�κ��� ���� ���� ���
                sound_timer <= SOUND_DURATION;  // Ÿ�̸� ����
            end
            
            // [Track 2 ����?]
            if (i_hit_t2 && i_btn_play[1]) begin
                o_judge <= 2'b11;        // Perfect!
                o_play_en <= 1;          // �Ҹ� ON
                o_cnt_limit <= i_curr_pitch_t2;  // LCD�κ��� ���� ���� ���
                sound_timer <= SOUND_DURATION;  // Ÿ�̸� ����
            end
            
            // ====================================================
            // 2. ���� �ʱ�ȭ (Auto Reset)
            // ====================================================
            else begin
                // 1ms ƽ�� ���� ������ ���� ���¸� �ʱ�ȭ�մϴ�.
                // (�̷��� �� �ϸ� Perfect�� ������ ������ �� ����)
                if (i_tick) begin
                    o_judge <= 0;       // IDLE ���·� ����
  
                    // �Ҹ� �ڵ� ���� ����
                    if (sound_timer > 0) begin
                        sound_timer <= sound_timer - 1;
                    end else begin
                        o_play_en <= 0; // �ð��� �� �Ǹ� �Ҹ� ����
                    end
                end
            end
        end
    end

endmodule