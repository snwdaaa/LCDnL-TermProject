module u_game_full_color_led (
    input clk,              // �ý��� Ŭ��
    input rst,              // ����
    input i_tick,           // 1ms ƽ (�ִϸ��̼� �ӵ� ������)
    input i_game_over,      // 1: ���� ����(�ִϸ��̼� ���), 0: ���� ��(���� ���)
    input [1:0] i_judge,    // ���� ��� (00:None, 01:Miss, 10:Normal, 11:Perfect)
    
    // ���� ��� �� (�� 4��Ʈ)
    output reg [3:0] o_fcl_r, // Red
    output reg [3:0] o_fcl_g, // Green
    output reg [3:0] o_fcl_b  // Blue
);

    // [1] ���� ���� (4��Ʈ��, ��� 1�̸� �ִ� ���) 
    // Red: R=1, G=0, B=0
    // Green: R=0, G=1, B=0
    // Yellow: R=1, G=1, B=0 (���� ȥ��)
    localparam COLOR_OFF = 12'h000;
    localparam COLOR_RED = 12'hF00;   // Miss
    localparam COLOR_YEL = 12'hFF0;   // Normal
    localparam COLOR_GRN = 12'h0F0;   // Perfect

    // [2] ���� ���� �ִϸ��̼� Ÿ�̸�
    reg [31:0] anim_cnt;
    reg [1:0] anim_step; // 0:Red -> 1:Yellow -> 2:Green ���� ����
    parameter ANIM_SPEED = 500; // 500ms���� �� ����

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            anim_cnt <= 0;
            anim_step <= 0;
        end else if (i_game_over && i_tick) begin
            // ���� ���� ������ ���� Ÿ�̸� ����
            if (anim_cnt >= ANIM_SPEED - 1) begin
                anim_cnt <= 0;
                // 0 -> 1 -> 2 -> 0 ... ���� �ݺ� (�Ǵ� ���߰� ���� ����)
                if (anim_step >= 2) anim_step <= 0;
                else anim_step <= anim_step + 1;
            end else begin
                anim_cnt <= anim_cnt + 1;
            end
        end
    end

    // [3] ��� ���� (�켱���� MUX)
    // Combinational Logic: �Է� ���¿� ���� ��� ���� ����
    always @(*) begin
        if (rst) begin
            {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_OFF;
        end 
        else if (i_game_over) begin
            // [��� 1] ���� ����: ���� �ִϸ��̼� ���
            case (anim_step)
                0: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_RED;
                1: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_YEL;
                2: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_GRN;
                default: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_OFF;
            endcase
        end 
        else begin
            // [��� 2] ���� ��: ���� ��� ���
            case (i_judge)
                2'b01: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_RED; // Miss
                2'b10: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_YEL; // Normal
                2'b11: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_GRN; // Perfect
                default: {o_fcl_r, o_fcl_g, o_fcl_b} = COLOR_OFF; // ��� ����
            endcase
        end
    end

endmodule