// ��Ʈ ������
// ���� ���� �ð��� ���� �Ǻ� ������ ���� ��ȣ ����

module note_gen (
    input clk,
    input rst,
    input [31:0] i_cur_time, // game_timer���� ���� ���� �ð� (ms)
    
    output reg o_note_t1,    // Track 1 (����) ��Ʈ ���� ��ȣ (1ƽ ���� 1)
    output reg o_note_t2,    // Track 2 (�Ʒ���) ��Ʈ ���� ��ȣ
    output reg [31:0] o_gen_pitch, // ������ ��Ʈ�� ���ļ� ��
    output reg o_game_end    // �뷡�� �������� �˸��� ��ȣ
);

    // ==========================================
    // �Ǻ� ������ �ϵ��ڵ�
    // ==========================================
    
    reg [31:0] note_time [0:NOTE_COUNT-1]; // �ð� ����
    reg [1:0]  note_track [0:NOTE_COUNT-1]; // Ʈ�� ���� (1:����, 2:�Ʒ���, 3:����)
    reg [31:0] note_pitch [0:NOTE_COUNT-1]; // ���� ���� �迭

// ==========================================
    // ? Smoke on the Water (Intro Riff)
    // ==========================================
    
    // 1. ���ļ� ��� ���� (50MHz Ŭ�� ���� ī���� ��)
    // ����: 50,000,000 / (���ļ� * 2)
    localparam G3  = 127551; // �� (196 Hz)
    localparam Bb3 = 107296; // ��b (233 Hz)
    localparam C4  = 95556;  // �� (262 Hz)
    localparam Db4 = 90197;  // ��b (277 Hz) - 6�� ����

    // ��Ʈ ���� (�� 12�� ��Ʈ�� ������ ����)
    parameter NOTE_COUNT = 12;
    
    reg [31:0] note_time  [0:NOTE_COUNT-1];
    reg [1:0]  note_track [0:NOTE_COUNT-1];
    reg [31:0] note_pitch [0:NOTE_COUNT-1];

    initial begin
        // BPM 112 ����: 4����ǥ(1��) ? 536ms, 8����ǥ(�ݹ�) ? 268ms
        // ���� �ð�: 1000ms (1�� ��� �� ����)

        // --- [Part 1] 0 - 3 - 5 ---
        note_time[0] = 1000;       note_track[0] = 2; note_pitch[0] = G3;  // �Ʒ���
        note_time[1] = 1536;       note_track[1] = 1; note_pitch[1] = Bb3; // ����
        note_time[2] = 2072;       note_track[2] = 2; note_pitch[2] = C4;  // �Ʒ���

        // --- [Part 2] 0 - 3 - 6 - 5 --- 
        // (���Ⱑ 5��, 6�� ��Ʈ �����Դϴ�!)
        note_time[3] = 3144;       note_track[3] = 1; note_pitch[3] = G3;  // ����
        note_time[4] = 3680;       note_track[4] = 2; note_pitch[4] = Bb3; // �Ʒ���
        
        // [����] 5��, 6���� ��ġ�� �ʰ� Ȯ���� �и�!
        note_time[5] = 4216;       note_track[5] = 1; note_pitch[5] = Db4; // ���� ("��")
        note_time[6] = 4752;       note_track[6] = 2; note_pitch[6] = C4;  // �Ʒ��� ("��~")

        // --- [Part 3] 0 - 3 - 5 - 3 - 0 ---
        note_time[7] = 5556;       note_track[7] = 1; note_pitch[7] = G3;  // ����
        note_time[8] = 6092;       note_track[8] = 2; note_pitch[8] = Bb3; // �Ʒ���
        note_time[9] = 6628;       note_track[9] = 1; note_pitch[9] = C4;  // ����
        note_time[10] = 7164;      note_track[10] = 2; note_pitch[10] = Bb3; // �Ʒ���
        note_time[11] = 7700;      note_track[11] = 1; note_pitch[11] = G3;  // ����
    end

    // ==========================================
    // ������ ���� (FSM)
    // ==========================================
    reg [31:0] note_idx; // ���� �� ��° ��Ʈ�� ��ٸ��� ������ (������)

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            note_idx <= 0;
            o_note_t1 <= 0;
            o_note_t2 <= 0;
            o_gen_pitch <= 0;
            o_game_end <= 0;
        end else begin
            o_note_t1 <= 0;
            o_note_t2 <= 0;

            // �뷡�� ���� �� �����ٸ�
            if (note_idx < NOTE_COUNT) begin
                // ���� �ð��� ��Ʈ�� �ð��� ���ų� ��������? (������ ��� ��� >= ���)
                if (i_cur_time >= note_time[note_idx]) begin
                    // ���� ���� ���
                    o_gen_pitch <= note_pitch[note_idx];
                    
                    // �ش� Ʈ���� ��ȣ �߻�
                    if (note_track[note_idx] == 1) 
                        o_note_t1 <= 1;
                    
                    if (note_track[note_idx] == 2) 
                        o_note_t2 <= 1;

                    // ���� ��Ʈ�� ������ �̵�
                    note_idx <= note_idx + 1;
                end
            end else begin
                // ��� ��Ʈ�� �� �������� ���� ���� ��ȣ
                // (������ ��Ʈ ������ ���� �ڿ� ������ ������ ���⼭ �ð� üũ�� �� �ص� ��)
                o_game_end <= 1;
            end
        end
    end

endmodule